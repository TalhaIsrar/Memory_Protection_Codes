module hamming_sec_decoder(
    input  [20:0] in_code;
    output [15:0] out_data;
    output error_corrected;
);

    always @(*) begin
        

    end
endmodule