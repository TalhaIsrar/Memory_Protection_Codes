module hamming_sec_encoder(
    input  [15:0] input_data;
    output [20:0] output_code;
);

    always @(*) begin
        

    end
endmodule