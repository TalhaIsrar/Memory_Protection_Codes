module hamming_sec_decoder(
    input  [11:0] in_code;
    output [7:0] out_data;
    output error_corrected;
);


endmodule